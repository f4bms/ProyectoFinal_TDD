module extend(
    input logic [23:0] Instruction,
    input logic [1:0] ImmSrc, // 00: Sign Extend, 01: Zero Extend, 10: PC Relative, 11: Unused
    output logic [31:0] ExtImm // Extensión de Instrucción
);

    always_comb begin
        case (ImmSrc)
            2'b00: ExtImm = {24'b0, Instruction[7:0]}; 
            2'b01: ExtImm = {20'b0, Instruction[11:0]}; 
            2'b10: ExtImm = {{6{Instruction[23]}}, Instruction[23:0], 2'b00};
            2'b11: ExtImm = 32'b0; // No se usa, pero se define para completar el caso
            default: ExtImm = 32'b0; // Manejo de caso por defecto
        endcase
    end
endmodule