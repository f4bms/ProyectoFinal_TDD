module sprites(
	output logic [3:0] door_open [0:17471],
	output logic [3:0] door_closed [0:17471],
	output logic [3:0] heart [0:439],
	output logic [3:0] player_1[0:719],
	output logic [3:0] player_2[0:719]
	);

logic [3:0] p1 [0:719] = '{
4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0100,
 4'b0100,
 4'b0100,
 4'b0100,
 4'b0100,
 4'b0100,
 4'b0100,
 4'b0100,
 4'b0100,
 4'b0100,
 4'b0100,
 4'b0100,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0100,
 4'b0100,
 4'b0100,
 4'b0100,
 4'b0100,
 4'b0100,
 4'b0100,
 4'b0100,
 4'b0100,
 4'b0100,
 4'b0100,
 4'b0100,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0100,
 4'b0100,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0100,
 4'b0100,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0100,
 4'b0100,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0100,
 4'b0100,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0111,
 4'b0111,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0111,
 4'b0111,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0111,
 4'b0111,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0111,
 4'b0111,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0111,
 4'b0111,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0111,
 4'b0111,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b1000,
 4'b1000,
 4'b1000,
 4'b1000,
 4'b1000,
 4'b1000,
 4'b1000,
 4'b1000,
 4'b1000,
 4'b1000,
 4'b1000,
 4'b1000,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b1000,
 4'b1000,
 4'b1000,
 4'b1000,
 4'b1000,
 4'b1000,
 4'b1000,
 4'b1000,
 4'b1000,
 4'b1000,
 4'b1000,
 4'b1000,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0111,
 4'b0111,
 4'b1000,
 4'b1000,
 4'b1000,
 4'b1000,
 4'b1000,
 4'b1000,
 4'b1000,
 4'b1000,
 4'b0111,
 4'b0111,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0111,
 4'b0111,
 4'b1000,
 4'b1000,
 4'b1000,
 4'b1000,
 4'b1000,
 4'b1000,
 4'b1000,
 4'b1000,
 4'b0111,
 4'b0111,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0100,
 4'b0100,
 4'b0100,
 4'b0100,
 4'b0111,
 4'b0111,
 4'b1000,
 4'b1000,
 4'b1000,
 4'b1000,
 4'b1000,
 4'b1000,
 4'b1000,
 4'b1000,
 4'b0111,
 4'b0111,
 4'b0100,
 4'b0100,
 4'b0100,
 4'b0100,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0100,
 4'b0100,
 4'b0100,
 4'b0100,
 4'b0111,
 4'b0111,
 4'b1000,
 4'b1000,
 4'b1000,
 4'b1000,
 4'b1000,
 4'b1000,
 4'b1000,
 4'b1000,
 4'b0111,
 4'b0111,
 4'b0100,
 4'b0100,
 4'b0100,
 4'b0100,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0100,
 4'b0100,
 4'b0100,
 4'b0100,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0100,
 4'b0100,
 4'b0100,
 4'b0100,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0100,
 4'b0100,
 4'b0100,
 4'b0100,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0100,
 4'b0100,
 4'b0100,
 4'b0100,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110
};

assign player_1 = p1;

logic [3:0] p2 [0:719] = '{
4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0100,
 4'b0100,
 4'b0100,
 4'b0100,
 4'b0100,
 4'b0100,
 4'b0100,
 4'b0100,
 4'b0100,
 4'b0100,
 4'b0100,
 4'b0100,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0100,
 4'b0100,
 4'b0100,
 4'b0100,
 4'b0100,
 4'b0100,
 4'b0100,
 4'b0100,
 4'b0100,
 4'b0100,
 4'b0100,
 4'b0100,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0100,
 4'b0100,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0100,
 4'b0100,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0100,
 4'b0100,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0100,
 4'b0100,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0111,
 4'b0111,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0111,
 4'b0111,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0111,
 4'b0111,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0111,
 4'b0111,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0111,
 4'b0111,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0111,
 4'b0111,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b1100,
 4'b1100,
 4'b1100,
 4'b1100,
 4'b1100,
 4'b1100,
 4'b1100,
 4'b1100,
 4'b1100,
 4'b1100,
 4'b1100,
 4'b1100,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b1100,
 4'b1100,
 4'b1100,
 4'b1100,
 4'b1100,
 4'b1100,
 4'b1100,
 4'b1100,
 4'b1100,
 4'b1100,
 4'b1100,
 4'b1100,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0111,
 4'b0111,
 4'b1100,
 4'b1100,
 4'b1100,
 4'b1100,
 4'b1100,
 4'b1100,
 4'b1100,
 4'b1100,
 4'b0111,
 4'b0111,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0111,
 4'b0111,
 4'b1100,
 4'b1100,
 4'b1100,
 4'b1100,
 4'b1100,
 4'b1100,
 4'b1100,
 4'b1100,
 4'b0111,
 4'b0111,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0100,
 4'b0100,
 4'b0100,
 4'b0100,
 4'b0111,
 4'b0111,
 4'b1100,
 4'b1100,
 4'b1100,
 4'b1100,
 4'b1100,
 4'b1100,
 4'b1100,
 4'b1100,
 4'b0111,
 4'b0111,
 4'b0100,
 4'b0100,
 4'b0100,
 4'b0100,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0100,
 4'b0100,
 4'b0100,
 4'b0100,
 4'b0111,
 4'b0111,
 4'b1100,
 4'b1100,
 4'b1100,
 4'b1100,
 4'b1100,
 4'b1100,
 4'b1100,
 4'b1100,
 4'b0111,
 4'b0111,
 4'b0100,
 4'b0100,
 4'b0100,
 4'b0100,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0100,
 4'b0100,
 4'b0100,
 4'b0100,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0100,
 4'b0100,
 4'b0100,
 4'b0100,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0100,
 4'b0100,
 4'b0100,
 4'b0100,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0100,
 4'b0100,
 4'b0100,
 4'b0100,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110
};

assign player_2 = p2;

logic [3:0] closed [0:17471] = '{
4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0110,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0010,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0110,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0110,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1010,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0110,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0110,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b1010,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1101,
 4'b1010,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1101,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0111,
 4'b0111,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1101,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b1001,
 4'b1001,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b1001,
 4'b1001,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0110,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b1001,
 4'b1001,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b1001,
 4'b1001,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b1001,
 4'b1001,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1101,
 4'b1010,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0111,
 4'b0111,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0111,
 4'b0111,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1010,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1010,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1010,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1010,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b0100,
 4'b0100,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b0100,
 4'b0100,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b0100,
 4'b0100,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b0100,
 4'b0100,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b0100,
 4'b0100,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b0100,
 4'b0100,
 4'b0100,
 4'b0100,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b0100,
 4'b0100,
 4'b0100,
 4'b0100,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b0100,
 4'b0100,
 4'b0100,
 4'b0100,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b0100,
 4'b0100,
 4'b0100,
 4'b0100,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b0100,
 4'b0100,
 4'b0100,
 4'b0100,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b0100,
 4'b0100,
 4'b0100,
 4'b0100,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b0100,
 4'b0100,
 4'b0100,
 4'b0100,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b0100,
 4'b0100,
 4'b0100,
 4'b0100,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b0100,
 4'b0100,
 4'b0100,
 4'b0100,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b0100,
 4'b0100,
 4'b0100,
 4'b0100,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b0100,
 4'b0100,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b0100,
 4'b0100,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b0100,
 4'b0100,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b0100,
 4'b0100,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b0100,
 4'b0100,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0110,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1101,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0111,
 4'b0111,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0111,
 4'b0111,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1010,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b0110,
 4'b0101,
 4'b0110,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b0110,
 4'b0110,
 4'b0110,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b0110,
 4'b0110,
 4'b0100,
 4'b0100,
 4'b0100,
 4'b0110,
 4'b0110,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1010,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b0110,
 4'b0110,
 4'b0110,
 4'b0110,
 4'b0100,
 4'b0110,
 4'b0110,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b0110,
 4'b0110,
 4'b0100,
 4'b0100,
 4'b0100,
 4'b0110,
 4'b0110,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b0110,
 4'b0110,
 4'b0100,
 4'b0100,
 4'b0100,
 4'b0011,
 4'b0110,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b0110,
 4'b0110,
 4'b0100,
 4'b0100,
 4'b0100,
 4'b0110,
 4'b0110,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1101,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0111,
 4'b0111,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b0110,
 4'b0110,
 4'b0100,
 4'b0100,
 4'b0100,
 4'b0110,
 4'b0110,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1010,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b0110,
 4'b0110,
 4'b0110,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b0100,
 4'b0110,
 4'b0110,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0111,
 4'b0111,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b0100,
 4'b0100,
 4'b0110,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1010,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b0100,
 4'b0100,
 4'b0110,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1010,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b0100,
 4'b0110,
 4'b0110,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1010,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b0110,
 4'b0100,
 4'b0110,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1010,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b0110,
 4'b0110,
 4'b0110,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b0100,
 4'b0110,
 4'b0110,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b0110,
 4'b0110,
 4'b0110,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b0110,
 4'b0110,
 4'b0110,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1010,
 4'b1101,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b0110,
 4'b0110,
 4'b0110,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b0011,
 4'b0110,
 4'b0110,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0111,
 4'b0111,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b0110,
 4'b0110,
 4'b0110,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b0110,
 4'b0101,
 4'b0110,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b0101,
 4'b0011,
 4'b0110,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b0100,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0111,
 4'b0111,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b0011,
 4'b0110,
 4'b0100,
 4'b0100,
 4'b0100,
 4'b0100,
 4'b0110,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b0110,
 4'b0110,
 4'b0100,
 4'b0100,
 4'b0100,
 4'b0110,
 4'b0110,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b0110,
 4'b0110,
 4'b0100,
 4'b0100,
 4'b0100,
 4'b0110,
 4'b0101,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1101,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b0110,
 4'b0110,
 4'b0110,
 4'b0100,
 4'b0100,
 4'b0110,
 4'b0110,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1010,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b0110,
 4'b0110,
 4'b0100,
 4'b0100,
 4'b0100,
 4'b0110,
 4'b0110,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0110,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b0110,
 4'b0110,
 4'b0110,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b0110,
 4'b0110,
 4'b0110,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b1001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b1001,
 4'b0111,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0111,
 4'b0111,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b1001,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0111,
 4'b0111,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b1001,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1010,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1010,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1010,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1010,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b0100,
 4'b0100,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b0100,
 4'b0100,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b0100,
 4'b0100,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b0100,
 4'b0100,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b0100,
 4'b0100,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b0100,
 4'b0100,
 4'b0100,
 4'b0100,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b0100,
 4'b0100,
 4'b0100,
 4'b0100,
 4'b1010,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b0100,
 4'b0100,
 4'b0100,
 4'b0100,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b0100,
 4'b0100,
 4'b0100,
 4'b0100,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b0100,
 4'b0100,
 4'b0100,
 4'b0100,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b0100,
 4'b0100,
 4'b0100,
 4'b0100,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b0100,
 4'b0100,
 4'b0100,
 4'b0100,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b0100,
 4'b0100,
 4'b0100,
 4'b0100,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b0100,
 4'b0100,
 4'b0100,
 4'b0100,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b0100,
 4'b0100,
 4'b0100,
 4'b0100,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b1010,
 4'b0100,
 4'b0100,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b0100,
 4'b0100,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b1010,
 4'b0100,
 4'b0100,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b0100,
 4'b0100,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b0100,
 4'b0100,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0110,
 4'b0011,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0101,
 4'b0111,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b1001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b1001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0111,
 4'b0111,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0111,
 4'b0111,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1101,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110
};
 
assign door_closed = closed;

logic [3:0] open [0:17471] = '{
4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0110,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0010,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0110,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0110,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0110,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0110,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0110,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0110,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0110,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b1001,
 4'b1001,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b1001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b1001,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b1001,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b1001,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0110,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b1001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b1001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110
};

assign door_open = open;

logic [3:0] heart_mem [0:439] = '{
4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b1111,
 4'b1111,
 4'b1111,
 4'b1111,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b1111,
 4'b1111,
 4'b1111,
 4'b1111,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b1111,
 4'b1111,
 4'b0000,
 4'b0000,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b1111,
 4'b1111,
 4'b1111,
 4'b1111,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b1111,
 4'b1111,
 4'b1111,
 4'b1111,
 4'b0000,
 4'b0000,
 4'b1111,
 4'b1111,
 4'b0111,
 4'b0111,
 4'b1111,
 4'b1111,
 4'b1111,
 4'b1111,
 4'b1111,
 4'b1111,
 4'b1111,
 4'b1111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b1111,
 4'b1111,
 4'b0000,
 4'b0000,
 4'b1111,
 4'b1111,
 4'b1111,
 4'b1111,
 4'b0111,
 4'b0111,
 4'b1111,
 4'b1111,
 4'b1111,
 4'b1111,
 4'b1111,
 4'b1111,
 4'b1111,
 4'b1111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b1111,
 4'b1111,
 4'b0000,
 4'b0000,
 4'b1111,
 4'b1111,
 4'b1111,
 4'b1111,
 4'b1111,
 4'b1111,
 4'b1111,
 4'b1111,
 4'b1111,
 4'b1111,
 4'b1111,
 4'b1111,
 4'b1111,
 4'b1111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b1111,
 4'b1111,
 4'b1111,
 4'b1111,
 4'b1111,
 4'b1111,
 4'b1111,
 4'b1111,
 4'b1111,
 4'b1111,
 4'b1111,
 4'b1111,
 4'b1111,
 4'b1111,
 4'b1111,
 4'b1111,
 4'b1111,
 4'b1111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b1111,
 4'b1111,
 4'b1111,
 4'b1111,
 4'b1111,
 4'b1111,
 4'b1111,
 4'b1111,
 4'b1111,
 4'b1111,
 4'b1111,
 4'b1111,
 4'b1111,
 4'b1111,
 4'b1111,
 4'b1111,
 4'b1111,
 4'b1111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b1111,
 4'b1111,
 4'b1111,
 4'b1111,
 4'b1111,
 4'b1111,
 4'b1111,
 4'b1111,
 4'b1111,
 4'b1111,
 4'b1111,
 4'b1111,
 4'b1111,
 4'b1111,
 4'b1111,
 4'b1111,
 4'b1111,
 4'b1111,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b1111,
 4'b1111,
 4'b1111,
 4'b1111,
 4'b1111,
 4'b1111,
 4'b1111,
 4'b1111,
 4'b1111,
 4'b1111,
 4'b1111,
 4'b1111,
 4'b1111,
 4'b1111,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b1111,
 4'b1111,
 4'b1111,
 4'b1111,
 4'b1111,
 4'b1111,
 4'b1111,
 4'b1111,
 4'b1111,
 4'b1111,
 4'b1111,
 4'b1111,
 4'b1111,
 4'b1111,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b1111,
 4'b1111,
 4'b1111,
 4'b1111,
 4'b1111,
 4'b1111,
 4'b1111,
 4'b1111,
 4'b1111,
 4'b1111,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b1111,
 4'b1111,
 4'b1111,
 4'b1111,
 4'b1111,
 4'b1111,
 4'b1111,
 4'b1111,
 4'b1111,
 4'b1111,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b1111,
 4'b1111,
 4'b1111,
 4'b1111,
 4'b1111,
 4'b1111,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b1111,
 4'b1111,
 4'b1111,
 4'b1111,
 4'b1111,
 4'b1111,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b1111,
 4'b1111,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b1111,
 4'b1111,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110
};

assign heart = heart_mem;

endmodule