module sprites(
	output logic [23:0] door_open [0:20271],
	output logic [23:0] door_closed [0:17471]
	//output logic [23:0] heart [0:399]
	);

logic [23:0] memory [0:17471] = '{
4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0111,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0111,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0111,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0111,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0111,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0111,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0111,
 4'b0000,
 4'b0000,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0111,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0000,
 4'b0111,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0111,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0110,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0111,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0010,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0110,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0110,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0111,
 4'b0000,
 4'b0000,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1010,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0000,
 4'b0000,
 4'b0111,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0110,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0111,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0111,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0110,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0111,
 4'b0000,
 4'b0000,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b1010,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1101,
 4'b1010,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0111,
 4'b0111,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1101,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0000,
 4'b0111,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0111,
 4'b0111,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1101,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b1001,
 4'b1001,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b1001,
 4'b1001,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0110,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b1001,
 4'b1001,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0000,
 4'b0111,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b1001,
 4'b1001,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b1001,
 4'b1001,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1101,
 4'b1010,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0111,
 4'b0111,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0111,
 4'b0111,
 4'b0000,
 4'b0000,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b0111,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b0111,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b0111,
 4'b1010,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0111,
 4'b0111,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0111,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0001,
 4'b0111,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0111,
 4'b0001,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0111,
 4'b0111,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b0111,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b0111,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b1001,
 4'b1001,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1000,
 4'b1001,
 4'b1001,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b0111,
 4'b0111,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1010,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b0111,
 4'b1101,
 4'b1101,
 4'b1010,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1010,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b0111,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1010,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1000,
 4'b1001,
 4'b1001,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b0100,
 4'b0100,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b0100,
 4'b0100,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b0100,
 4'b0100,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b0100,
 4'b0100,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b0100,
 4'b0100,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1000,
 4'b1001,
 4'b1001,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b0100,
 4'b0100,
 4'b0100,
 4'b0100,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b0100,
 4'b0100,
 4'b0100,
 4'b0100,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b0100,
 4'b0100,
 4'b0100,
 4'b0100,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b0100,
 4'b0100,
 4'b0100,
 4'b0100,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b0100,
 4'b0100,
 4'b0100,
 4'b0100,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1000,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b0100,
 4'b0100,
 4'b0100,
 4'b0100,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b0100,
 4'b0100,
 4'b0100,
 4'b0100,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b0100,
 4'b0100,
 4'b0100,
 4'b0100,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b0100,
 4'b0100,
 4'b0100,
 4'b0100,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b0111,
 4'b0111,
 4'b1011,
 4'b0100,
 4'b0100,
 4'b0100,
 4'b0100,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1000,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0001,
 4'b0111,
 4'b0001,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b0100,
 4'b0100,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b0111,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b0100,
 4'b0100,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b0100,
 4'b0100,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b0100,
 4'b0100,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b0100,
 4'b0100,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1000,
 4'b1001,
 4'b1001,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b0111,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b0111,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1000,
 4'b1001,
 4'b1001,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0110,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1000,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0111,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b1000,
 4'b1000,
 4'b1000,
 4'b1000,
 4'b1000,
 4'b1000,
 4'b1000,
 4'b1000,
 4'b1000,
 4'b1000,
 4'b1000,
 4'b1000,
 4'b1000,
 4'b1000,
 4'b1000,
 4'b1000,
 4'b1000,
 4'b1000,
 4'b1000,
 4'b1000,
 4'b1000,
 4'b1000,
 4'b1000,
 4'b1000,
 4'b1000,
 4'b1000,
 4'b1000,
 4'b1000,
 4'b1000,
 4'b1000,
 4'b1000,
 4'b1000,
 4'b1000,
 4'b1000,
 4'b1000,
 4'b1000,
 4'b1000,
 4'b1000,
 4'b1000,
 4'b1000,
 4'b1000,
 4'b1000,
 4'b1000,
 4'b1000,
 4'b1000,
 4'b1000,
 4'b1000,
 4'b1000,
 4'b1000,
 4'b1000,
 4'b1000,
 4'b1000,
 4'b1000,
 4'b1000,
 4'b1000,
 4'b1000,
 4'b1000,
 4'b1000,
 4'b1000,
 4'b1000,
 4'b1000,
 4'b1000,
 4'b1000,
 4'b1000,
 4'b1000,
 4'b1000,
 4'b1000,
 4'b1000,
 4'b1000,
 4'b1000,
 4'b1000,
 4'b1000,
 4'b1000,
 4'b1000,
 4'b1000,
 4'b1000,
 4'b1000,
 4'b1000,
 4'b1000,
 4'b1000,
 4'b1000,
 4'b1000,
 4'b1000,
 4'b1000,
 4'b1000,
 4'b1000,
 4'b1000,
 4'b1001,
 4'b1001,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0111,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b0111,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1101,
 4'b1010,
 4'b0111,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0111,
 4'b0111,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b0111,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b0111,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b0111,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b0111,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b0111,
 4'b1101,
 4'b0111,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0111,
 4'b0111,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b0111,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b0111,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b0111,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1010,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b0111,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b0110,
 4'b0111,
 4'b0110,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b0111,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b0110,
 4'b0110,
 4'b0110,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b0111,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b0110,
 4'b0110,
 4'b0100,
 4'b0100,
 4'b0100,
 4'b0110,
 4'b0110,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1010,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b0110,
 4'b0110,
 4'b0111,
 4'b0111,
 4'b0100,
 4'b0110,
 4'b0110,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b0111,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b0110,
 4'b0110,
 4'b0100,
 4'b0100,
 4'b0100,
 4'b0110,
 4'b0110,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b0111,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b0110,
 4'b0110,
 4'b0100,
 4'b0100,
 4'b0100,
 4'b0111,
 4'b0110,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b0110,
 4'b0110,
 4'b0100,
 4'b0100,
 4'b0100,
 4'b0110,
 4'b0110,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1101,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0111,
 4'b0111,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b0110,
 4'b0110,
 4'b0100,
 4'b0100,
 4'b0100,
 4'b0110,
 4'b0110,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1010,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b0110,
 4'b0110,
 4'b0110,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b0111,
 4'b0110,
 4'b0110,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b0111,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0111,
 4'b0111,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b0111,
 4'b0111,
 4'b0110,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1010,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b0111,
 4'b0111,
 4'b0110,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1010,
 4'b1011,
 4'b0111,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1010,
 4'b0111,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0111,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b0111,
 4'b0110,
 4'b0110,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1010,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b0110,
 4'b0111,
 4'b0110,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b0111,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1010,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b0111,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b0110,
 4'b0110,
 4'b0110,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b0111,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b0111,
 4'b1011,
 4'b0111,
 4'b0110,
 4'b0110,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b0111,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b0110,
 4'b0110,
 4'b0110,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b0110,
 4'b0110,
 4'b0110,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1010,
 4'b1101,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0111,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b0110,
 4'b0110,
 4'b0110,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b0111,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b0111,
 4'b0110,
 4'b0110,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b0111,
 4'b1010,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0111,
 4'b0111,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b0110,
 4'b0110,
 4'b0110,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b0111,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b0110,
 4'b0111,
 4'b0110,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b0111,
 4'b0111,
 4'b0110,
 4'b1011,
 4'b0111,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b0111,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b0111,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b0111,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0111,
 4'b0111,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b0111,
 4'b0110,
 4'b0111,
 4'b0100,
 4'b0100,
 4'b0111,
 4'b0110,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b0110,
 4'b0110,
 4'b0100,
 4'b0100,
 4'b0100,
 4'b0110,
 4'b0110,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b0110,
 4'b0110,
 4'b0100,
 4'b0100,
 4'b0100,
 4'b0110,
 4'b0111,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1101,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b0110,
 4'b0110,
 4'b0111,
 4'b0111,
 4'b0100,
 4'b0110,
 4'b0110,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1010,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b0111,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b0110,
 4'b0110,
 4'b0100,
 4'b0100,
 4'b0100,
 4'b0110,
 4'b0111,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b0111,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0110,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b0110,
 4'b0110,
 4'b0110,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b0111,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b0110,
 4'b0110,
 4'b0110,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b0111,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b0111,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b0111,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0111,
 4'b0111,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0111,
 4'b0111,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b1000,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1000,
 4'b1001,
 4'b1001,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b1000,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1010,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1010,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1010,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1010,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1000,
 4'b1001,
 4'b1001,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0111,
 4'b0001,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b1000,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b0100,
 4'b0100,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b0100,
 4'b0100,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b0100,
 4'b0100,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b0100,
 4'b0100,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b0100,
 4'b0100,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1000,
 4'b1001,
 4'b1001,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b1000,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b0100,
 4'b0100,
 4'b0100,
 4'b0100,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b0100,
 4'b0111,
 4'b0100,
 4'b0100,
 4'b1010,
 4'b1011,
 4'b0111,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b0111,
 4'b1011,
 4'b0100,
 4'b0100,
 4'b0100,
 4'b0100,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b0100,
 4'b0100,
 4'b0100,
 4'b0100,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b0100,
 4'b0100,
 4'b0100,
 4'b0100,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1000,
 4'b1001,
 4'b1001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b1000,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b0111,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b0100,
 4'b0100,
 4'b0100,
 4'b0100,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b0100,
 4'b0111,
 4'b0100,
 4'b0100,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b0100,
 4'b0100,
 4'b0100,
 4'b0100,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b0100,
 4'b0100,
 4'b0100,
 4'b0100,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b0100,
 4'b0100,
 4'b0100,
 4'b0100,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1000,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b1000,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b0111,
 4'b0100,
 4'b0100,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b0100,
 4'b0100,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b0100,
 4'b0100,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b0100,
 4'b0100,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b0100,
 4'b0100,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1000,
 4'b1001,
 4'b1001,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b1000,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1000,
 4'b1001,
 4'b1001,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0110,
 4'b0011,
 4'b1000,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1000,
 4'b1001,
 4'b1001,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b1000,
 4'b1001,
 4'b1001,
 4'b1000,
 4'b1000,
 4'b1000,
 4'b1000,
 4'b1000,
 4'b1000,
 4'b1000,
 4'b1000,
 4'b1000,
 4'b1000,
 4'b1000,
 4'b1000,
 4'b1000,
 4'b1000,
 4'b1000,
 4'b1000,
 4'b1000,
 4'b1000,
 4'b1000,
 4'b1000,
 4'b1000,
 4'b1000,
 4'b1000,
 4'b1000,
 4'b1000,
 4'b1000,
 4'b1000,
 4'b1000,
 4'b1000,
 4'b1000,
 4'b1000,
 4'b1000,
 4'b1000,
 4'b1000,
 4'b1000,
 4'b1000,
 4'b1000,
 4'b1000,
 4'b1000,
 4'b1000,
 4'b1000,
 4'b1000,
 4'b1000,
 4'b1000,
 4'b1000,
 4'b1000,
 4'b1000,
 4'b1000,
 4'b1000,
 4'b1000,
 4'b1000,
 4'b1000,
 4'b1000,
 4'b1000,
 4'b1000,
 4'b1000,
 4'b1000,
 4'b1000,
 4'b1000,
 4'b1000,
 4'b1000,
 4'b1000,
 4'b1000,
 4'b1000,
 4'b1000,
 4'b1000,
 4'b1000,
 4'b1000,
 4'b1000,
 4'b1000,
 4'b1000,
 4'b1000,
 4'b1000,
 4'b1000,
 4'b1000,
 4'b1000,
 4'b1000,
 4'b1000,
 4'b1000,
 4'b1000,
 4'b1000,
 4'b1000,
 4'b1000,
 4'b1000,
 4'b1000,
 4'b1000,
 4'b1001,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0111,
 4'b0111,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0111,
 4'b0111,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1101,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0000,
 4'b0000,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0000,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0000, 
 4'b0000
};
 
assign door_closed = memory;

logic [23:0] open [0:20271] = '{
4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1010,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b0111,
 4'b1100,
 4'b1100,
 4'b1100,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1010,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b0111,
 4'b1100,
 4'b1100,
 4'b1100,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1010,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b0111,
 4'b1100,
 4'b1100,
 4'b1100,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1010,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b0111,
 4'b1100,
 4'b1100,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1010,
 4'b1101,
 4'b0111,
 4'b1101,
 4'b1101,
 4'b0111,
 4'b1100,
 4'b1100,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0011,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1010,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b0111,
 4'b1100,
 4'b1100,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b0111,
 4'b1100,
 4'b1100,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0011,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b0111,
 4'b1101,
 4'b0111,
 4'b0111,
 4'b1100,
 4'b1100,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0011,
 4'b0011,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1010,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b0111,
 4'b0111,
 4'b1100,
 4'b1100,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0011,
 4'b0011,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1010,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b0111,
 4'b1101,
 4'b1101,
 4'b0111,
 4'b1100,
 4'b1100,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0011,
 4'b0011,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1010,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b0111,
 4'b1101,
 4'b1101,
 4'b0111,
 4'b1100,
 4'b1100,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1010,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b0111,
 4'b1100,
 4'b1100,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1010,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b0111,
 4'b1100,
 4'b1100,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b0111,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1010,
 4'b0111,
 4'b1101,
 4'b0111,
 4'b1101,
 4'b0111,
 4'b1100,
 4'b1100,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b0111,
 4'b0111,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1010,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b0111,
 4'b1100,
 4'b1100,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b0111,
 4'b0111,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1010,
 4'b0111,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b0111,
 4'b1100,
 4'b1100,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1010,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b0111,
 4'b1100,
 4'b1100,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1010,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b0111,
 4'b1100,
 4'b1100,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1010,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b0111,
 4'b1100,
 4'b1100,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b0010,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1010,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b0111,
 4'b1100,
 4'b1100,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b0011,
 4'b0011,
 4'b0001,
 4'b0111,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1010,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b0111,
 4'b1100,
 4'b1100,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b0011,
 4'b0011,
 4'b0001,
 4'b0111,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1010,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b0111,
 4'b1100,
 4'b1100,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b1001,
 4'b0111,
 4'b1001,
 4'b1010,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b0111,
 4'b1100,
 4'b1100,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1010,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b0111,
 4'b1100,
 4'b1100,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1010,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b0111,
 4'b1100,
 4'b1100,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1010,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b0111,
 4'b1100,
 4'b1100,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1010,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b0111,
 4'b1100,
 4'b1100,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0111,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1010,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b0111,
 4'b1100,
 4'b1100,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0101,
 4'b0101,
 4'b0111,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1010,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b0111,
 4'b1100,
 4'b1100,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1010,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b0111,
 4'b1100,
 4'b1100,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b0111,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1010,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b0111,
 4'b1100,
 4'b1100,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b0111,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1010,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b0111,
 4'b1100,
 4'b1100,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b0111,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b0111,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b1001,
 4'b0111,
 4'b1001,
 4'b1010,
 4'b1101,
 4'b1101,
 4'b0111,
 4'b0111,
 4'b1101,
 4'b1101,
 4'b0111,
 4'b1100,
 4'b1100,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b0111,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b0111,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1010,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b0111,
 4'b1100,
 4'b1100,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b0111,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b0111,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b1001,
 4'b1001,
 4'b1010,
 4'b1101,
 4'b1101,
 4'b0111,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b0111,
 4'b1100,
 4'b0111,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b0111,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1001,
 4'b0111,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b0111,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b1001,
 4'b1001,
 4'b1010,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b0111,
 4'b1100,
 4'b1100,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b0111,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1001,
 4'b0111,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b0111,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b1001,
 4'b1001,
 4'b1010,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b0111,
 4'b1100,
 4'b1100,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b0111,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1001,
 4'b0111,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b0111,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b0111,
 4'b1001,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0111,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0111,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b1001,
 4'b1001,
 4'b1010,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b0111,
 4'b1100,
 4'b1100,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b0111,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b0111,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0111,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0111,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b1001,
 4'b1001,
 4'b1010,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b0111,
 4'b1100,
 4'b1100,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b0111,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b1001,
 4'b1001,
 4'b1010,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b0111,
 4'b1100,
 4'b1100,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b0111,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b1001,
 4'b1001,
 4'b1010,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b0111,
 4'b1100,
 4'b1100,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b0111,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b1001,
 4'b1001,
 4'b1010,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b0111,
 4'b1100,
 4'b1100,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b0111,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b1001,
 4'b1001,
 4'b1010,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b0111,
 4'b1100,
 4'b1100,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b0111,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b1001,
 4'b1001,
 4'b1010,
 4'b1101,
 4'b1101,
 4'b0111,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b0111,
 4'b1100,
 4'b1100,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b0111,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b1001,
 4'b1001,
 4'b1010,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b0111,
 4'b1100,
 4'b1100,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b0111,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b1001,
 4'b1001,
 4'b1010,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b0111,
 4'b1100,
 4'b1100,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b0111,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b1001,
 4'b1001,
 4'b1010,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b0111,
 4'b1100,
 4'b1100,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b1001,
 4'b1001,
 4'b1010,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0111,
 4'b0111,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b1001,
 4'b1001,
 4'b1010,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b0111,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b1001,
 4'b1001,
 4'b1010,
 4'b1101,
 4'b1101,
 4'b1001,
 4'b1001,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b0111,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b1001,
 4'b1001,
 4'b1010,
 4'b1101,
 4'b1101,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b0111,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0111,
 4'b0111,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b1001,
 4'b1001,
 4'b1010,
 4'b1101,
 4'b1101,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b0111,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b1001,
 4'b1001,
 4'b1010,
 4'b1101,
 4'b1101,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b0111,
 4'b0111,
 4'b1011,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b0111,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b1001,
 4'b1001,
 4'b1010,
 4'b1101,
 4'b1101,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b0111,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b1001,
 4'b1001,
 4'b1010,
 4'b1101,
 4'b1101,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b0100,
 4'b0100,
 4'b0100,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b0111,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b1001,
 4'b1001,
 4'b1010,
 4'b1101,
 4'b1101,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b0111,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b0100,
 4'b0100,
 4'b0100,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b0101,
 4'b0111,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b1001,
 4'b1001,
 4'b1010,
 4'b1101,
 4'b1101,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b0100,
 4'b0100,
 4'b0100,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b0100,
 4'b0100,
 4'b0100,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b0101,
 4'b0111,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b1001,
 4'b1001,
 4'b1010,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b0100,
 4'b0100,
 4'b0100,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b0101,
 4'b0111,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b1001,
 4'b1001,
 4'b1010,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b0100,
 4'b0100,
 4'b0100,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b0100,
 4'b0100,
 4'b0100,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b0101,
 4'b0111,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b1001,
 4'b1001,
 4'b1010,
 4'b1101,
 4'b0111,
 4'b1101,
 4'b1101,
 4'b0111,
 4'b1101,
 4'b1101,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b0100,
 4'b0100,
 4'b0100,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b0101,
 4'b0111,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0111,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b1001,
 4'b1001,
 4'b1010,
 4'b0111,
 4'b0111,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b0100,
 4'b0100,
 4'b0100,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0111,
 4'b0111,
 4'b0101,
 4'b0111,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0111,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b1001,
 4'b1001,
 4'b1010,
 4'b0111,
 4'b0111,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b0100,
 4'b0100,
 4'b0100,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1001,
 4'b1001,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0101,
 4'b0111,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0111,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b1001,
 4'b1001,
 4'b1010,
 4'b0111,
 4'b0111,
 4'b1101,
 4'b1101,
 4'b0111,
 4'b1101,
 4'b0111,
 4'b1100,
 4'b1100,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b0100,
 4'b0100,
 4'b0100,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1001,
 4'b1001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b1001,
 4'b1001,
 4'b1010,
 4'b0111,
 4'b0111,
 4'b1101,
 4'b1101,
 4'b0111,
 4'b1101,
 4'b0111,
 4'b1100,
 4'b1100,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b0100,
 4'b0100,
 4'b0100,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1001,
 4'b1001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0111,
 4'b0111,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b1001,
 4'b1001,
 4'b1010,
 4'b0111,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b1100,
 4'b1100,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b0100,
 4'b0100,
 4'b0100,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b0101,
 4'b0111,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b1001,
 4'b1001,
 4'b1010,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b0111,
 4'b0111,
 4'b1100,
 4'b1100,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b0111,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b0100,
 4'b0100,
 4'b0100,
 4'b1011,
 4'b0111,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b0101,
 4'b0111,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b1001,
 4'b1001,
 4'b1010,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b0111,
 4'b1100,
 4'b1100,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b0111,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b0100,
 4'b0100,
 4'b0100,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b0101,
 4'b0111,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b1001,
 4'b1001,
 4'b1010,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b0111,
 4'b1100,
 4'b1100,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b0111,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b0101,
 4'b0111,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b1001,
 4'b1001,
 4'b1010,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b0111,
 4'b1100,
 4'b1100,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b0111,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b0101,
 4'b0111,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b1001,
 4'b1001,
 4'b1010,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b0111,
 4'b1100,
 4'b1100,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b0111,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b0101,
 4'b0111,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b1001,
 4'b1001,
 4'b1010,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b0111,
 4'b1100,
 4'b1100,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b0111,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b0101,
 4'b0111,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b1001,
 4'b1001,
 4'b1010,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b0111,
 4'b1100,
 4'b1100,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b0111,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b0111,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b1001,
 4'b1001,
 4'b1010,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b0111,
 4'b1100,
 4'b1100,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b0111,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b1001,
 4'b1001,
 4'b1010,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b0111,
 4'b1101,
 4'b1101,
 4'b0111,
 4'b1100,
 4'b1100,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b0111,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b0111,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0111,
 4'b0111,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b1001,
 4'b1001,
 4'b1010,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b0111,
 4'b1101,
 4'b1101,
 4'b0111,
 4'b1100,
 4'b1100,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b0111,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b0111,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0111,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b1001,
 4'b1001,
 4'b1010,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b0111,
 4'b1100,
 4'b1100,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b0111,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b0111,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0111,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b1001,
 4'b1001,
 4'b1010,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b0111,
 4'b1100,
 4'b1100,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b0111,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0111,
 4'b0111,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0111,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b1001,
 4'b1001,
 4'b1010,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b0111,
 4'b1100,
 4'b1100,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b0111,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b0111,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0001,
 4'b0111,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0111,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b1001,
 4'b1001,
 4'b1010,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b0111,
 4'b1100,
 4'b1100,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b0110,
 4'b0110,
 4'b0110,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b0111,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b0111,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0111,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0111,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b1001,
 4'b1001,
 4'b1010,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b0111,
 4'b1100,
 4'b1100,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b0110,
 4'b0110,
 4'b0110,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b0111,
 4'b1001,
 4'b1101,
 4'b0111,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b0111,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b0111,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0111,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0111,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b1001,
 4'b1001,
 4'b1010,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b0111,
 4'b1100,
 4'b1100,
 4'b1011,
 4'b0110,
 4'b0110,
 4'b0100,
 4'b0100,
 4'b0100,
 4'b0110,
 4'b0110,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b0111,
 4'b1001,
 4'b1101,
 4'b0111,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b0111,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b0111,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0111,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b1001,
 4'b1001,
 4'b1010,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b0111,
 4'b1100,
 4'b1100,
 4'b1011,
 4'b0111,
 4'b0110,
 4'b0100,
 4'b0100,
 4'b0100,
 4'b0111,
 4'b0110,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b0111,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b0111,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b0111,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0111,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b1001,
 4'b1001,
 4'b1010,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b0111,
 4'b1100,
 4'b1100,
 4'b1011,
 4'b0111,
 4'b0110,
 4'b0100,
 4'b0100,
 4'b0100,
 4'b0111,
 4'b0110,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b0111,
 4'b1001,
 4'b1101,
 4'b0111,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b0111,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b0111,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0111,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b1001,
 4'b1001,
 4'b1010,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b0111,
 4'b1100,
 4'b1100,
 4'b1011,
 4'b0111,
 4'b0110,
 4'b0100,
 4'b0100,
 4'b0100,
 4'b0111,
 4'b0110,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b0111,
 4'b1001,
 4'b1101,
 4'b0111,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b0111,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b0111,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0111,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b1001,
 4'b1001,
 4'b1010,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b0111,
 4'b1101,
 4'b1101,
 4'b0111,
 4'b1100,
 4'b1100,
 4'b1011,
 4'b0111,
 4'b0110,
 4'b0100,
 4'b0100,
 4'b0100,
 4'b0111,
 4'b0110,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b0111,
 4'b1001,
 4'b1101,
 4'b0111,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b0111,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b0111,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b0111,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0111,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b1001,
 4'b1001,
 4'b1010,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b0111,
 4'b1100,
 4'b1100,
 4'b1011,
 4'b0110,
 4'b0110,
 4'b0100,
 4'b0100,
 4'b0100,
 4'b0111,
 4'b0110,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b0111,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b0111,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0111,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b1001,
 4'b1001,
 4'b1010,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b0111,
 4'b1100,
 4'b1100,
 4'b1011,
 4'b0110,
 4'b0110,
 4'b0100,
 4'b0100,
 4'b0100,
 4'b0110,
 4'b0110,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b0111,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b0111,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0111,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0111,
 4'b0111,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b1001,
 4'b1001,
 4'b1010,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b0111,
 4'b1100,
 4'b1100,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b0110,
 4'b0110,
 4'b0110,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b0111,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b0111,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b1001,
 4'b1001,
 4'b1010,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b0111,
 4'b1100,
 4'b1100,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b0110,
 4'b0110,
 4'b0110,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b0111,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b0111,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b0111,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b1001,
 4'b1001,
 4'b1010,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b0111,
 4'b1100,
 4'b1100,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b0110,
 4'b0111,
 4'b0110,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b0111,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b0111,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0111,
 4'b0111,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b1001,
 4'b1001,
 4'b1010,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b0111,
 4'b1100,
 4'b1100,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b0110,
 4'b0111,
 4'b0110,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b0111,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b0111,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b1001,
 4'b1001,
 4'b1010,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b0111,
 4'b1100,
 4'b1100,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b0110,
 4'b0111,
 4'b0110,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b0111,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b0111,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b1001,
 4'b1001,
 4'b1010,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b0111,
 4'b1100,
 4'b1100,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b0110,
 4'b0111,
 4'b0110,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b0111,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b0111,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b1001,
 4'b1001,
 4'b1010,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b0111,
 4'b1101,
 4'b1101,
 4'b0111,
 4'b1100,
 4'b1100,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b0110,
 4'b0111,
 4'b0110,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b0111,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b1001,
 4'b1001,
 4'b1010,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b0111,
 4'b1101,
 4'b1101,
 4'b0111,
 4'b1100,
 4'b1100,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b0110,
 4'b0111,
 4'b0110,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b0111,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b0111,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b1001,
 4'b1001,
 4'b1010,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b0111,
 4'b1100,
 4'b1100,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b0110,
 4'b0111,
 4'b0110,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b0111,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b0111,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b0111,
 4'b1001,
 4'b1101,
 4'b0111,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b1001,
 4'b1001,
 4'b1010,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b0111,
 4'b1100,
 4'b1100,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b0110,
 4'b0111,
 4'b0110,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b0111,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b0111,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b0111,
 4'b1001,
 4'b1101,
 4'b0111,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b1001,
 4'b1001,
 4'b1010,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b0111,
 4'b1100,
 4'b1100,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b0110,
 4'b0111,
 4'b0110,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b0111,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b0111,
 4'b1001,
 4'b1101,
 4'b0111,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b0111,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b0111,
 4'b1001,
 4'b1101,
 4'b0111,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b1001,
 4'b1001,
 4'b1010,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b0111,
 4'b1100,
 4'b1100,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b0110,
 4'b0111,
 4'b0110,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b0111,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b0111,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b0111,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b0111,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0111,
 4'b0111,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b1001,
 4'b1001,
 4'b1010,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b0111,
 4'b1100,
 4'b1100,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b0110,
 4'b0111,
 4'b0110,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b0111,
 4'b1001,
 4'b1101,
 4'b0111,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b0111,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0111,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b1001,
 4'b1001,
 4'b1010,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b0111,
 4'b1100,
 4'b1100,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b0110,
 4'b0111,
 4'b0110,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b0111,
 4'b1001,
 4'b1101,
 4'b0111,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b0111,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0111,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b1001,
 4'b1001,
 4'b1010,
 4'b1101,
 4'b0111,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b0111,
 4'b1100,
 4'b1100,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b0110,
 4'b0111,
 4'b0110,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b0111,
 4'b1001,
 4'b1101,
 4'b0111,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b0111,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0111,
 4'b0111,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0111,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b1001,
 4'b1001,
 4'b1010,
 4'b1101,
 4'b0111,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b0111,
 4'b1100,
 4'b1100,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b0110,
 4'b0111,
 4'b0110,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b0111,
 4'b1001,
 4'b1101,
 4'b0111,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b0111,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0111,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b1001,
 4'b1001,
 4'b1010,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b0111,
 4'b1100,
 4'b1100,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b0110,
 4'b0111,
 4'b0110,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b0111,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0111,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b1001,
 4'b1001,
 4'b1010,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b0111,
 4'b1100,
 4'b1100,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b0110,
 4'b0110,
 4'b0110,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b0111,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b0111,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0111,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0111,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0111,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b1001,
 4'b1001,
 4'b1010,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b0111,
 4'b1100,
 4'b1100,
 4'b1011,
 4'b0110,
 4'b0110,
 4'b0100,
 4'b0100,
 4'b0100,
 4'b0110,
 4'b0110,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b0111,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b0111,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0111,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0111,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b1001,
 4'b1001,
 4'b1010,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b0111,
 4'b1100,
 4'b1100,
 4'b1011,
 4'b0110,
 4'b0110,
 4'b0100,
 4'b0100,
 4'b0100,
 4'b0110,
 4'b0110,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b0111,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b0111,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b1001,
 4'b1001,
 4'b1010,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b0111,
 4'b1100,
 4'b1100,
 4'b1011,
 4'b0110,
 4'b0110,
 4'b0100,
 4'b0100,
 4'b0100,
 4'b0110,
 4'b0110,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b0111,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b1001,
 4'b1001,
 4'b1010,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b0111,
 4'b1100,
 4'b1100,
 4'b1011,
 4'b0110,
 4'b0110,
 4'b0100,
 4'b0100,
 4'b0100,
 4'b0110,
 4'b0110,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b1001,
 4'b1001,
 4'b1010,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b0111,
 4'b1100,
 4'b1100,
 4'b1011,
 4'b0110,
 4'b0110,
 4'b0100,
 4'b0100,
 4'b0100,
 4'b0110,
 4'b0110,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b0111,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b1001,
 4'b1001,
 4'b1010,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b0111,
 4'b1100,
 4'b1100,
 4'b1011,
 4'b0110,
 4'b0110,
 4'b0100,
 4'b0100,
 4'b0100,
 4'b0110,
 4'b0110,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b0111,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b1001,
 4'b1001,
 4'b1010,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b0111,
 4'b1100,
 4'b1100,
 4'b1011,
 4'b0110,
 4'b0110,
 4'b0100,
 4'b0100,
 4'b0100,
 4'b0110,
 4'b0110,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b0111,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0111,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0111,
 4'b0111,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b1001,
 4'b1001,
 4'b1010,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b0111,
 4'b1100,
 4'b1100,
 4'b1011,
 4'b0110,
 4'b0110,
 4'b0100,
 4'b0100,
 4'b0100,
 4'b0110,
 4'b0110,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b0111,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b1001,
 4'b1001,
 4'b1010,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b0111,
 4'b1100,
 4'b1100,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b0110,
 4'b0110,
 4'b0110,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b0111,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b1001,
 4'b1001,
 4'b1010,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b0111,
 4'b1100,
 4'b1100,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b0110,
 4'b0110,
 4'b0110,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b0111,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b0111,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0111,
 4'b0111,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b1001,
 4'b1001,
 4'b1010,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b0111,
 4'b1100,
 4'b1100,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b0111,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b1001,
 4'b1001,
 4'b1010,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b0111,
 4'b1100,
 4'b1100,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b1001,
 4'b1001,
 4'b1010,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b0111,
 4'b1100,
 4'b1100,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b0111,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b0111,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b1001,
 4'b1001,
 4'b1010,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b0111,
 4'b1100,
 4'b1100,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b1001,
 4'b1001,
 4'b1010,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b0111,
 4'b1100,
 4'b1100,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b1001,
 4'b1001,
 4'b1010,
 4'b0111,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b0111,
 4'b1100,
 4'b1100,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b1001,
 4'b1001,
 4'b1010,
 4'b1101,
 4'b1101,
 4'b0111,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b0111,
 4'b1100,
 4'b1100,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b0011,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b1001,
 4'b1001,
 4'b1010,
 4'b1101,
 4'b1101,
 4'b0111,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b0111,
 4'b1100,
 4'b1100,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b1001,
 4'b1001,
 4'b1010,
 4'b1101,
 4'b1101,
 4'b0111,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b0111,
 4'b1100,
 4'b1100,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b1001,
 4'b1001,
 4'b1010,
 4'b1101,
 4'b1101,
 4'b0111,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b0111,
 4'b1100,
 4'b1100,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0111,
 4'b0111,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b1001,
 4'b1001,
 4'b1010,
 4'b1101,
 4'b1101,
 4'b0111,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b0111,
 4'b1100,
 4'b1100,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0111,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b1001,
 4'b1001,
 4'b1010,
 4'b0111,
 4'b1101,
 4'b0111,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b0111,
 4'b1100,
 4'b1100,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b1001,
 4'b1001,
 4'b1010,
 4'b0111,
 4'b1101,
 4'b0111,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b0111,
 4'b1100,
 4'b1100,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0111,
 4'b0111,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0111,
 4'b0111,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b1001,
 4'b1001,
 4'b1010,
 4'b0111,
 4'b1101,
 4'b0111,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b0111,
 4'b1100,
 4'b1100,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b0100,
 4'b0100,
 4'b0100,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0111,
 4'b0111,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b1001,
 4'b1001,
 4'b1010,
 4'b0111,
 4'b1101,
 4'b0111,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b0111,
 4'b1100,
 4'b1100,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b0100,
 4'b0100,
 4'b0100,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0111,
 4'b0111,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b1001,
 4'b1001,
 4'b1010,
 4'b1101,
 4'b1101,
 4'b0111,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b0111,
 4'b1100,
 4'b1100,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b0100,
 4'b0100,
 4'b0100,
 4'b1011,
 4'b0111,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b0100,
 4'b0100,
 4'b0100,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0111,
 4'b0111,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b1001,
 4'b1001,
 4'b1010,
 4'b1101,
 4'b1101,
 4'b0111,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b0111,
 4'b1100,
 4'b1100,
 4'b1011,
 4'b0111,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b0100,
 4'b0100,
 4'b0100,
 4'b1011,
 4'b0111,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0111,
 4'b0111,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b1001,
 4'b1001,
 4'b1010,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b0111,
 4'b1100,
 4'b1100,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b0111,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b0100,
 4'b0100,
 4'b0100,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0111,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b1001,
 4'b1001,
 4'b1010,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b0100,
 4'b0100,
 4'b0100,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0111,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b1001,
 4'b1001,
 4'b1010,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b0100,
 4'b0100,
 4'b0100,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0111,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b1001,
 4'b1001,
 4'b1010,
 4'b1101,
 4'b1101,
 4'b1001,
 4'b1001,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1010,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b0100,
 4'b0100,
 4'b0100,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b0100,
 4'b0100,
 4'b0100,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0111,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b1001,
 4'b1001,
 4'b1010,
 4'b1101,
 4'b1101,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b0100,
 4'b0100,
 4'b0100,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0111,
 4'b0111,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0111,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b1001,
 4'b1001,
 4'b1010,
 4'b1101,
 4'b1101,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b0100,
 4'b0100,
 4'b0100,
 4'b1011,
 4'b1011,
 4'b0111,
 4'b0111,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0111,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b1001,
 4'b1001,
 4'b1010,
 4'b1101,
 4'b1101,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b0100,
 4'b0100,
 4'b0100,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0111,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b1001,
 4'b1001,
 4'b1010,
 4'b1101,
 4'b1101,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b0100,
 4'b0100,
 4'b0100,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0111,
 4'b0111,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0111,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b1001,
 4'b1001,
 4'b1010,
 4'b1101,
 4'b1101,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b0100,
 4'b0100,
 4'b0100,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0111,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b1001,
 4'b1001,
 4'b1010,
 4'b1101,
 4'b1101,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0111,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b1001,
 4'b1001,
 4'b1010,
 4'b1101,
 4'b1101,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0111,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b1001,
 4'b1001,
 4'b1010,
 4'b1101,
 4'b1101,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0111,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b1001,
 4'b1001,
 4'b1010,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1010,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0111,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b1001,
 4'b1001,
 4'b1010,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0111,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b1001,
 4'b1001,
 4'b1010,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b0111,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b1001,
 4'b1001,
 4'b1010,
 4'b1101,
 4'b0111,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b0111,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b1001,
 4'b1001,
 4'b1010,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b0111,
 4'b1100,
 4'b1100,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b1001,
 4'b1001,
 4'b1010,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b0111,
 4'b1100,
 4'b1100,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b0111,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0010,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0111,
 4'b0111,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b0101,
 4'b1001,
 4'b1001,
 4'b1010,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b0111,
 4'b1100,
 4'b1100,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b0111,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0011,
 4'b0010,
 4'b0001,
 4'b0001,
 4'b0001,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b1001,
 4'b1001,
 4'b1010,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b0111,
 4'b1100,
 4'b1100,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b0111,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b1001,
 4'b1001,
 4'b1010,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b0111,
 4'b1100,
 4'b1100,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b0111,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b0111,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1001,
 4'b1001,
 4'b1010,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b0111,
 4'b1100,
 4'b1100,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b0111,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1001,
 4'b1001,
 4'b1010,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b0111,
 4'b1100,
 4'b1100,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b0111,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1001,
 4'b1001,
 4'b1010,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b0111,
 4'b1100,
 4'b1100,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b0111,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1001,
 4'b1001,
 4'b1010,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b0111,
 4'b1100,
 4'b1100,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1001,
 4'b1001,
 4'b1010,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b0111,
 4'b1100,
 4'b1100,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b0111,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1001,
 4'b1001,
 4'b1010,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b0111,
 4'b1100,
 4'b1100,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1001,
 4'b1001,
 4'b1010,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b0111,
 4'b1100,
 4'b1100,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1001,
 4'b1001,
 4'b1010,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b0111,
 4'b1100,
 4'b1100,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b0111,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1001,
 4'b1001,
 4'b1010,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b0111,
 4'b1101,
 4'b0111,
 4'b1100,
 4'b1100,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1001,
 4'b1001,
 4'b1010,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b0111,
 4'b1100,
 4'b1100,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1001,
 4'b1001,
 4'b1010,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b0111,
 4'b1100,
 4'b1100,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1010,
 4'b1010,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1001,
 4'b1001,
 4'b1010,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b0111,
 4'b1100,
 4'b1100,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1001,
 4'b1001,
 4'b1010,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b0111,
 4'b1100,
 4'b1100,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1001,
 4'b1001,
 4'b1010,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b0111,
 4'b1100,
 4'b1100,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1001,
 4'b1001,
 4'b1010,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b0111,
 4'b1100,
 4'b1100,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1001,
 4'b1001,
 4'b1010,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b0111,
 4'b1100,
 4'b1100,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1001,
 4'b1001,
 4'b1010,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b0111,
 4'b1100,
 4'b1100,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1001,
 4'b1001,
 4'b1010,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b0111,
 4'b1100,
 4'b1100,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1101,
 4'b1101,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1001,
 4'b1001,
 4'b1010,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b0111,
 4'b1100,
 4'b1100,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1001,
 4'b1001,
 4'b1010,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b0111,
 4'b1100,
 4'b1100,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b0111,
 4'b1001,
 4'b1001,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1001,
 4'b1001,
 4'b1010,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b0111,
 4'b1100,
 4'b1100,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1001,
 4'b1001,
 4'b1010,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b0111,
 4'b1100,
 4'b1100,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1001,
 4'b1001,
 4'b1010,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b0111,
 4'b1100,
 4'b1100,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1001,
 4'b1001,
 4'b1010,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b1101,
 4'b0111,
 4'b1100,
 4'b1100,
 4'b1011,
 4'b1011,
 4'b1011,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1001,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110,
 4'b1110
};

assign door_open = open;

endmodule